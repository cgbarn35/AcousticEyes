`timescale 100ns / 10ps


`define HalfClockPeriod 1.6

module PDMTest;

initial begin 
	$dumpfile("out.vcd");
	$dumpvars;
end

//INPUT
reg CLK;
reg RST;
reg [3000:0] testData; //TODO VERIFIY TEST LENGTH
reg [11:0] cnt;
reg sftData;
//OUTPUT
wire CLKDIV;
wire [15:0] OUT;

ClockDivider C0(//TODO PARAMETERIZE CLOCK DIVISION
	CLK,
	RST,
	CLKDIV
	);

	CICNR16 #(3) uut (
		.clk(CLK),
		.clkdiv(CLKDIV),
		.rst(RST),
		.x_in(sftData),
		.y_out(OUT)
		);


		initial begin 
			CLK = 0;
			RST = 0;
			cnt = 0;
			testData = 'b110101010101010101010101011010101010110101010110101011010110101101011010110101101011011011010110110110110101101101101101110110110110110111011011011101110110111011101101110111011101110111101110111011110111101111011101111101111011110111110111110111110111110111111011111101111111011111101111111101111111101111111110111111111101111111111101111111111111011111111111111101111111111111111111101111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111110111111111111111111111111110111111111111111111101111111111111101111111111111011111111111011111111101111111110111111110111111101111111011111101111110111111011111011111011111011111011110111101111011110111101111011101111011101110111011101110111011101110110111011101101101110110110111011011011011011011011011011011010110110110101101011011010110101101011010101101010110101011010101010110101010101010101101010101010101010100101010101010101001010101010010101001010100101010010100101001010010100100101001001001010010010010010010010010010010010010001001001000100100010010001000100100010001000100010000100010001000010001000010000100001000010000010000100000100000100000100000010000001000000100000001000000010000000010000000010000000000100000000001000000000000100000000000000010000000000000000001000000000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000100000000000000001000000000000010000000000001000000000010000000001000000001000000010000000100000001000000100000010000010000010000010000010000010000100001000010000100001000100001000100010001000100010001000100010001001000100100010010010001001001001001001001001001001001001001001010010010100100101001010010100101001010100101010010101001010101010010101010101010101010101001101010101010101010101010110101010101101010110101011010101101011010110101101011011010110110110101101101101101101101101101101101101101110110111011011011101110110111011101110111011101110111011110111011110111101110111110111101111011111011110111110111110111111011111101111110111111011111111011111110111111110111111111101111111111011111111111101111111111111011111111111111111011111111111111111111110111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111110111111111111111111111110111111111111111110111111111111110111111111110111111111110111111111011111111011111111011111110111111101111110111111011111011111101111101111011111011110111101111011110111101111011101110111101110111011101110111011101101110111011011011101101110110110;
			#100
			RST = 1;
			#100
			RST = 0;

			#10000 //TODO DETERMINE
			$finish;
	end

	always begin                                                 
		#`HalfClockPeriod CLK = ~CLK;                         
	end

	always @(posedge CLK or posedge RST) begin                                                 
		if(RST) begin 
			cnt = 0;
			sftData = 0;
		end
		else begin
		cnt = cnt + 1;
		sftData = testData[cnt];
	end
end

	endmodule

	module ClockDivider(
		input clk,
		input rst,
		output reg clkdiv
		);
		parameter N = 16;

		reg[6:0] cnt;
		initial begin 
			cnt = 0;
			clkdiv = 0;
		end


		always @(posedge clk) begin 
			if(rst) begin 
				cnt = 0;
				clkdiv = 0;
			end
			cnt <= cnt + 1;
			if(cnt >= N-1) begin
				cnt <= 0;
				clkdiv <= ~clkdiv;
			end
		end
		endmodule
